/*
 Copyright 2013 Ray Salemi

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at

 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 */
module top;
import tinyalu_pkg::*;
`include "tinyalu_macros.svh"

tinyalu DUT (.A(bfm.A), .B(bfm.B), .op(bfm.op),
    .clk(bfm.clk), .reset_n(bfm.reset_n),
    .start(bfm.start), .done(bfm.done), .result(bfm.result));

tinyalu_bfm bfm();

testbench testbench_h;


initial begin
    testbench_h = new(bfm);
    testbench_h.execute();
end

endmodule : top


